module common

import time

pub const (
	max_page_limit = 10
	sleep_duration = time.millisecond * 400
)
