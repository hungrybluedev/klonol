module main

enum Provider {
	github
	gitea
}

enum Action {
	list
	clone
	pull
}
