module main

enum Action {
	list
	clone
	pull
}
