module main

enum Provider {
	github
	gitea
}
